danny is lame in STD_LOGIC
