braden is lame in STD_LOGIC
