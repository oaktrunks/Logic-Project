danny is cool in STD_LOGIC