library IEEE; use IEEE.STD_Logic_1164.all;
entity LogicProject is
port(instruction: in STD_LOGIC_VECTOR (15 downto 0);
EXE, UPD: in STD_LOGIC;
enADD, enXOR, enMOVREGTOREG, enMOVDATA, enINC, enDEC, enROL, enROR, enNEG, enOUT: out STD_LOGIC;
end;
architecture decoder of LogicProject is
begin
UPD <=
enADD <=
enXOR <=
enMOVREGTOREG <=
enMOVDATA <=
enINC <=
enDEC <=
enROL <=
enROR <=
enNEG <=
enOUT <=
end;
